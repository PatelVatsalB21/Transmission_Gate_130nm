* C:\Users\Vatsal\eSim-Workspace\CMOS_Transmission_Gate\CMOS_Transmission_Gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/28/2021 12:14:37 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  IN -CONTROL OUT IN mosfet_p		
M2  OUT CONTROL IN IN mosfet_n		
v2  -CONTROL GND pulse		
v1  IN GND pulse		
v3  CONTROL GND pulse		
U1  IN plot_v1		
U2  -CONTROL plot_v1		
U3  CONTROL plot_v1		
U4  OUT plot_v1		

.end
